library verilog;
use verilog.vl_types.all;
entity memoria_4x3_vlg_vec_tst is
end memoria_4x3_vlg_vec_tst;
