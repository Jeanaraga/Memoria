library verilog;
use verilog.vl_types.all;
entity memoria_4x3_vlg_check_tst is
    port(
        O0              : in     vl_logic;
        O1              : in     vl_logic;
        O2              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end memoria_4x3_vlg_check_tst;
